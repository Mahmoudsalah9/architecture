LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;