LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY Execute IS
    PORT (

        Clk : IN STD_LOGIC;
        Rst : IN STD_LOGIC;
        

    );
END ENTITY;

ARCHITECTURE Execute_Design OF Execute IS






BEGIN
END;