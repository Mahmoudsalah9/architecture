LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY Decode IS
    PORT (

        Clk : IN STD_LOGIC;
        Rst : IN STD_LOGIC;
        Data_After : IN STD_LOGIC;

    );
END ENTITY;

ARCHITECTURE Decode_Design OF Decode IS






BEGIN
END;